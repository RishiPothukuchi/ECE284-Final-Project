`timescale 1ns/1ps

module core_tb;

parameter bw = 4;
parameter psum_bw = 16;
parameter len_kij = 9;
parameter len_onij = 16;
parameter col = 8;
parameter row = 8;
parameter len_nij = 36;

// pruning param
parameter PRUNING_MODE = 0;  // 0: no prune 1: unstructured 2: structured
parameter SPARSITY = 50;     // For unstructured, % of weights to zero (0-100)
parameter PRUNE_LAYER = 3;   // For structured which kij layer to zero (0-8)

// pruning save
reg [31:0] pruned_wt;
integer zero_ct;
integer nibble_idx;
integer rando_val;

reg clk = 0;
reg reset = 1;

wire [34:0] inst_q; 

reg [1:0]  inst_w_q = 0; 
reg [bw*row-1:0] D_xmem_q = 0;
reg CEN_xmem = 1;
reg WEN_xmem = 1;
reg [10:0] A_xmem = 0;
reg CEN_xmem_q = 1;
reg WEN_xmem_q = 1;
reg [10:0] A_xmem_q = 0;
reg CEN_pmem = 1;
reg WEN_pmem = 1;
reg [10:0] A_pmem = 0;
reg CEN_pmem_q = 1;
reg WEN_pmem_q = 1;
reg [10:0] A_pmem_q = 0;
reg ofifo_rd_q = 0;
reg ififo_wr_q = 0;
reg ififo_rd_q = 0;
reg l0_rd_q = 0;
reg l0_wr_q = 0;
reg execute_q = 0;
reg load_q = 0;
reg acc_q = 0;
reg acc = 0;
reg bypass = 0;
reg bypass_q = 0;

reg [1:0]  inst_w; 
reg [bw*row-1:0] D_xmem;
reg [psum_bw*col-1:0] answer;


reg ofifo_rd;
reg ififo_wr;
reg ififo_rd;
reg l0_rd;
reg l0_wr;
reg execute;
reg load;
reg [8*30:1] stringvar;
reg [8*30:1] w_file_name;
wire ofifo_valid;
wire [col*psum_bw-1:0] sfp_out;

integer x_file, x_scan_file ; // file_handler
integer w_file, w_scan_file ; // file_handler
integer acc_file, acc_scan_file ; // file_handler
integer out_file, out_scan_file ; // file_handler
integer captured_data; 
integer t, i, j, k, kij;
integer error;

assign inst_q[34] = bypass_q;
assign inst_q[33] = acc_q;
assign inst_q[32] = CEN_pmem_q;
assign inst_q[31] = WEN_pmem_q;
assign inst_q[30:20] = A_pmem_q;
assign inst_q[19]   = CEN_xmem_q;
assign inst_q[18]   = WEN_xmem_q;
assign inst_q[17:7] = A_xmem_q;
assign inst_q[6]   = ofifo_rd_q;
assign inst_q[5]   = ififo_wr_q;
assign inst_q[4]   = ififo_rd_q;
assign inst_q[3]   = l0_rd_q;
assign inst_q[2]   = l0_wr_q;
assign inst_q[1]   = execute_q; 
assign inst_q[0]   = load_q; 


core  #(.bw(bw), .col(col), .row(row)) core_instance (
	.clk(clk), 
	.inst(inst_q),
	.ofifo_valid(ofifo_valid),
        .D_xmem(D_xmem_q), 
        .sfp_out(sfp_out), 
	.reset(reset)); 


initial begin 

  inst_w   = 0; 
  D_xmem   = 0;
  CEN_xmem = 1;
  WEN_xmem = 1;
  A_xmem   = 0;
  ofifo_rd = 0;
  ififo_wr = 0;
  ififo_rd = 0;
  l0_rd    = 0;
  l0_wr    = 0;
  execute  = 0;
  load     = 0;

  $dumpfile("core_tb.vcd");
  $dumpvars(0,core_tb);

  x_file = $fopen("activation_tile0.txt", "r");
  // Following three lines are to remove the first three comment lines of the file
  x_scan_file = $fscanf(x_file,"%s", captured_data);
  x_scan_file = $fscanf(x_file,"%s", captured_data);
  x_scan_file = $fscanf(x_file,"%s", captured_data);

  //////// Reset /////////
  #0.5 clk = 1'b0;   reset = 1;
  #0.5 clk = 1'b1; 

  for (i=0; i<10 ; i=i+1) begin
    #0.5 clk = 1'b0;
    #0.5 clk = 1'b1;  
  end

  #0.5 clk = 1'b0;   reset = 0;
  #0.5 clk = 1'b1; 

  #0.5 clk = 1'b0;   
  #0.5 clk = 1'b1;   
  /////////////////////////

  /////// Activation data writing to memory ///////
  for (t=0; t<len_nij; t=t+1) begin  
    #0.5 clk = 1'b0;  x_scan_file = $fscanf(x_file,"%32b", D_xmem); WEN_xmem = 0; CEN_xmem = 0; if (t>0) A_xmem = A_xmem + 1;
    #0.5 clk = 1'b1;   
  end

  #0.5 clk = 1'b0;  WEN_xmem = 1;  CEN_xmem = 1; A_xmem = 0;
  #0.5 clk = 1'b1; 

  $fclose(x_file);
  /////////////////////////////////////////////////


  for (kij=0; kij<9; kij=kij+1) begin  // kij loop

    case(kij)
     0: w_file_name = "weight_itile0_otile0_kij0.txt";
     1: w_file_name = "weight_itile0_otile0_kij1.txt";
     2: w_file_name = "weight_itile0_otile0_kij2.txt";
     3: w_file_name = "weight_itile0_otile0_kij3.txt";
     4: w_file_name = "weight_itile0_otile0_kij4.txt";
     5: w_file_name = "weight_itile0_otile0_kij5.txt";
     6: w_file_name = "weight_itile0_otile0_kij6.txt";
     7: w_file_name = "weight_itile0_otile0_kij7.txt";
     8: w_file_name = "weight_itile0_otile0_kij8.txt";
    endcase
    

    w_file = $fopen(w_file_name, "r");
    // Following three lines are to remove the first three comment lines of the file
    w_scan_file = $fscanf(w_file,"%s", captured_data);
    w_scan_file = $fscanf(w_file,"%s", captured_data);
    w_scan_file = $fscanf(w_file,"%s", captured_data);

    #0.5 clk = 1'b0;   reset = 1;
    #0.5 clk = 1'b1; 

    for (i=0; i<10 ; i=i+1) begin
      #0.5 clk = 1'b0;
      #0.5 clk = 1'b1;  
    end

    #0.5 clk = 1'b0;   reset = 0;
    #0.5 clk = 1'b1; 

    #0.5 clk = 1'b0;   
    #0.5 clk = 1'b1;   





    /////// Kernel data writing to memory ///////

    A_xmem = 11'b10000000000;


	if (PRUNING_MODE == 1) begin
        $display("kij=%d: Unstructured pruning, %d sparsity", kij, SPARSITY);
    end
    else if (PRUNING_MODE == 2 && kij == PRUNE_LAYER) begin
        $display("kij=%d: Structured pruning", kij);
    end
    else if (PRUNING_MODE == 2) begin
        $display("kij=%d: No pruning, structured for layer %d", kij, PRUNE_LAYER);
    end
    else begin
        $display("kij=%0d: No pruning done", kij);
    end

	zero_ct = 0; 

    for (t=0; t<col; t=t+1) begin  
      #0.5 clk = 1'b0;
      
      w_scan_file = $fscanf(w_file,"%32b", D_xmem);
      
      pruned_wt = D_xmem; 
      
      case (PRUNING_MODE)
        
        // Mode 1: Unstructured
        1: begin
          for (nibble_idx = 0; nibble_idx < 8; nibble_idx = nibble_idx + 1) begin
            rando_val = $random % 100;
            if (rando_val < 0) begin
              rando_val = -rando_val; 
            end

            if (random_val < SPARSITY) begin
              pruned_wt[nibble_idx*4 +: 4] = 4'b0000;
              zero_ct = zero_ct + 1;
            end
          end
        end
        
        // Mode 2: Structured
        2: begin
          if (kij == PRUNE_LAYER) begin
            pruned_wt = 32'b0;
            zero_ct = zero_ct + 8; 
          end
        end
        
        // Mode 0: No pruning done
        default: begin
          pruned_wt = D_xmem;
        end
        
      endcase
      
      D_xmem = pruned_wt;
      WEN_xmem = 0;
      CEN_xmem = 0;
      
      if (t>0) begin
        A_xmem = A_xmem + 1;
      end
      
      #0.5 clk = 1'b1;  
    end
    
    if (PRUNING_MODE != 0) begin
      $display("kij=%0d: Zeroed %0d out of %0d weights (%.1f%%)", kij, zero_count, col*8, (zero_count*100.0)/(col*8));
    end
    
    #0.5 clk = 1'b0;  WEN_xmem = 1;  CEN_xmem = 1; A_xmem = 0;
    #0.5 clk = 1'b1; 
    /////////////////////////////////////


    /////// Kernel data writing to L0 ///////
    // prime SRAM and delay by a cycle, wr first addr to sram
    #0.5 clk = 1'b0;
    CEN_xmem = 0; // turn on SRAM
    WEN_xmem = 1; // read out mode
    A_xmem = 11'b10000000000;
    l0_wr = 0;
    #0.5 clk = 1'b1; 

    for (t=0; t<col; t=t+1) begin
      #0.5 clk = 1'b0;
 
      l0_wr = 1;
   
      if (t<col-1) begin
        A_xmem = A_xmem + 1;
      end 

      #0.5 clk = 1'b1;
    end

    // // iteration v3
    // // load in 0x407
    // #0.5 clk = 1'b0;
    // l0_wr = 1;
    // CEN_xmem = 1; // turn off SRAM but get its last output
    // #0.5 clk = 1'b1;

    #0.5 clk = 1'b0;
    CEN_xmem = 1;
    l0_wr = 0;
    #0.5 clk = 1'b1;

    // itervation v2
    // // turn off L0
    // #0.5 clk = 1'b0;
    // l0_wr = 0;
    // CEN_xmem = 1;
    // WEN_xmem = 1;
    // #0.5 clk = 1'b1;

  //   for (t=0; t<col; t=t+1) begin
  //   	#0.5 clk = 1'b0 CEN_xmem = 0; WEN_xmem = 1; A_xmem = 11'b10000000000 + t[10:0]; l0_wr = 1;
	// #0.5 clk = 1'b1;
  //   end

  //   #0.5 clk = 1'b0; l0_wr = 0; CEN_xmem = 1; WEN_xmem = 1;
  //   #0.5 clk = 1'b1;
    /////////////////////////////////////



    /////// Kernel loading to PEs ///////
    for (t=0; t<col+row; t=t+1) begin
      #0.5 clk = 1'b0; load = 1; l0_rd = 1;
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0; load = 0; l0_rd = 0;
    #0.5 clk = 1'b1;
    /////////////////////////////////////
  


    ////// provide some intermission to clear up the kernel loading ///
    #0.5 clk = 1'b0;  load = 0; l0_rd = 0;
    #0.5 clk = 1'b1;  
  

    for (i=0; i<10 ; i=i+1) begin
      #0.5 clk = 1'b0;
      #0.5 clk = 1'b1;  
    end
    /////////////////////////////////////



    /////// Activation data writing to L0 ///////
    #0.5 clk = 1'b0;
    CEN_xmem = 0;
    WEN_xmem = 1;
    A_xmem = 11'b00000000000;
    l0_wr = 0;
    #0.5 clk = 1'b1;


    for (t=0; t < len_nij; t=t+1) begin
      #0.5 clk = 1'b0;

      l0_wr = 1;

      if (t < len_nij - 1) begin
        A_xmem = A_xmem + 1;
      end 
      else begin
        CEN_xmem = 1;
      end
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0;
    l0_wr = 0;
    CEN_xmem = 1;
    WEN_xmem = 1;
    #0.5 clk = 1'b1;

  //   for (t=0; t<len_nij; t=t+1) begin
  //   	#0.5 clk = 1'b0; CEN_xmem = 0; WEN_xmem = 1; l0_wr = 1;
	// #0.5 clk = 1'b1; A_xmem = A_xmem + 1;
  //   end

  //   #0.5 clk = 1'b0; l0_wr = 0; CEN_xmem = 1; WEN_xmem = 1;
  //   #0.5 clk = 1'b1;
    /////////////////////////////////////

  // #0.5 clk = 1'b0;
  // l0_rd = 1;
  // execute = 0;
  // #0.5 clk = 1'b1;

    /////// Execution /////// ~36 cycles
    for (t=0; t<row+col+len_nij; t=t+1) begin
    	#0.5 clk = 1'b0; execute = 1; l0_rd = 1;
	    #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0; execute = 0; l0_rd = 0;
    #0.5 clk = 1'b1;
    /////////////////////////////////////



  //   ////// OFIFO READ ////////
  //   Ideally, OFIFO should be read while execution, but we have enough ofifo
  //   depth so we can fetch out after execution.
  // read out to and accum in sfu 16 times
    // wait 1 clk cycle for valid out
    // #0.5 clk = 1'b0;
    // acc = 0;
    // ofifo_rd = 1;
    // #0.5 clk = 1'b1;
    $display("\n===== PMEM Storage =====");
    #0.5 clk = 1'b0;
    acc = 0;                  // don't accumulate yet
    ofifo_rd = 1;             // read next PSUM, output to psum_in for SFU
    // CEN_pmem = 0;             // enable PMEM
    // WEN_pmem = 0;             // enable write on PMEM
    A_pmem = kij * len_onij;  // get starting address (i.e. kij=0 -> 0, kij=1 -> 16, kij=2 -> 32, etc.)
    bypass = 1;               // avoid acc + ReLU, just store raw PSUM result
    #0.5 clk = 1'b1;
    t=0;
    while (t < len_onij) begin // 2 cycle delay
      #0.5 clk = 1'b0; 
      if (ofifo_valid) begin
        ofifo_rd = 1;   // acc = 1;
        CEN_pmem = 0;   // enable PMEM
        WEN_pmem = 0;   // enable write on PMEM
        if ( t > 0 ) A_pmem = A_pmem + 1;
        t = t + 1;
        if (ofifo_valid && CEN_pmem == 0) begin
        $display("[KIJ=%0d, t=%0d] Writing to PMEM[%0d], sfp_out=%h", 
                kij, t, A_pmem, sfp_out);
        end
      end
      else begin
        ofifo_rd = 0;
        CEN_pmem = 1;
        WEN_pmem = 1;
        // acc = 0;
      end
      #0.5 clk = 1'b1;
    end

    #0.5 clk = 1'b0;
    ofifo_rd = 0;
    acc = 0;
    CEN_pmem = 1;     // disable PMEM
    WEN_pmem = 1;     // disable write on PMEM
    bypass = 0;       // remove bypass signal
    #0.5 clk = 1'b1;

    /////////////////////////////////////

  end  // end of kij loop



  ////////// Accumulation /////////
  out_file = $fopen("out.txt", "r");  

  acc_file = $fopen("acc.txt", "r");


  // Following three lines are to remove the first three comment lines of the file
  out_scan_file = $fscanf(out_file,"%s", answer); 
  out_scan_file = $fscanf(out_file,"%s", answer); 
  out_scan_file = $fscanf(out_file,"%s", answer); 

  error = 0;


  // drive ofifo, sfu, alongside answer checking to not lose data
  $display("############ Verification Start during accumulation #############");



  for (i=0; i<len_onij; i=i+1) begin 
    // assert read accumulate
    wait(ofifo_valid);

    #0.5 clk = 1'b0;
    ofifo_rd = 1;
    acc = 1;
    #0.5 clk = 1'b1;
    //read in one vector per loop it
    #0.5 clk = 1'b0;
    ofifo_rd = 0;
    acc = 0;
    #0.5 clk = 1'b1;
    // // flush and relu
    // #0.5 clk = 1'b0;
    // acc = 0;
    // #0.5 clk = 1'b1;
    // wait + calc
    #0.5 clk = 1'b0; #0.5 clk = 1'b1;
    #0.5 clk = 1'b0; #0.5 clk = 1'b1;

    out_scan_file = $fscanf(out_file,"%128b", answer); // reading from out file to answer
    if (sfp_out == answer)
      $display("%2d-th output featuremap Data matched! :D", i); 
    else begin
      $display("%2d-th output featuremap Data ERROR!!", i); 
      $display("sfpout: %128b", sfp_out);
      $display("answer: %128b", answer);
      $display("sfpout: %d", sfp_out);
      $display("answer: %d", answer);
      error = 1;
    end

    // if (i>0) begin
    //  out_scan_file = $fscanf(out_file,"%128b", answer); // reading from out file to answer
    //    if (sfp_out == answer)
    //      $display("%2d-th output featuremap Data matched! :D", i); 
    //    else begin
    //      $display("%2d-th output featuremap Data ERROR!!", i); 
    //      $display("sfpout: %128b", sfp_out);
    //      $display("answer: %128b", answer);
    //      error = 1;
    //    end
    // end
   
 
    // #0.5 clk = 1'b0; reset = 1;
    // #0.5 clk = 1'b1;  
    // #0.5 clk = 1'b0; reset = 0; 
    // #0.5 clk = 1'b1;  

    // for (j=0; j<len_kij+1; j=j+1) begin 

    //   #0.5 clk = 1'b0;   
    //     if (j<len_kij) begin CEN_pmem = 0; WEN_pmem = 1; acc_scan_file = $fscanf(acc_file,"%11b", A_pmem); end
    //                    else  begin CEN_pmem = 1; WEN_pmem = 1; end

    //     if (j>0)  acc = 1;  
    //   #0.5 clk = 1'b1;   
    // end

    // #0.5 clk = 1'b0; acc = 0;
    // #0.5 clk = 1'b1; 
  end


  if (error == 0) begin
  	$display("############ No error detected ##############"); 
  	$display("########### Project Completed !! ############"); 

  end

  $fclose(acc_file);
  //////////////////////////////////

  for (t=0; t<10; t=t+1) begin  
    #0.5 clk = 1'b0;  
    #0.5 clk = 1'b1;  
  end

  #10 $finish;

end

always @ (posedge clk) begin
   inst_w_q   <= inst_w; 
   D_xmem_q   <= D_xmem;
   CEN_xmem_q <= CEN_xmem;
   WEN_xmem_q <= WEN_xmem;
   A_pmem_q   <= A_pmem;
   CEN_pmem_q <= CEN_pmem;
   WEN_pmem_q <= WEN_pmem;
   A_xmem_q   <= A_xmem;
   ofifo_rd_q <= ofifo_rd;
   acc_q      <= acc;
   ififo_wr_q <= ififo_wr;
   ififo_rd_q <= ififo_rd;
   l0_rd_q    <= l0_rd;
   l0_wr_q    <= l0_wr ;
   execute_q  <= execute;
   load_q     <= load;
   bypass_q   <= bypass;
end





endmodule




